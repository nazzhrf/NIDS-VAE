`timescale 1ns / 1ps

module sqrt16slices

(
    input wire clk,          
    input wire rst,
    input wire sqrt_en,          
    input wire signed [15:0] x, 
    output wire signed [15:0] y
);
    // Wire to observe value
    wire signed [15:0] m16_w;
    wire signed [15:0] c16_w;
    wire signed [31:0] mx32_w;
    wire signed [15:0] mx16_w;

    // Register to save temporary value
    reg [3:0] cntr_sqrt;
    reg signed [15:0] m16_reg;
    reg signed [15:0] c16_reg;
    reg signed [31:0] mx32_reg;
    reg signed [15:0] mx16_reg;
    reg signed [15:0] y_reg;
    
    

    // Choose value of gradient m based on input x value
    assign m16_w =  (x >= 16'sb000000_0000000000 && x < 16'sb000000_0010101011)  ? 16'sb000010_0111001100 : // m1 = 2.4495
                    (x >= 16'sb000000_0010101011 && x < 16'sb000000_0101010101)  ? 16'sb000001_0000001111 : // m2 = 1.0146
                    (x >= 16'sb000000_0101010101 && x < 16'sb000000_1000000000)  ? 16'sb000000_1100011101 : // m3 = 0.7785
                    (x >= 16'sb000000_1000000000 && x <= 16'sb000000_1010101011) ? 16'sb000000_1010100000 : // m4 = 0.6563
                    (x >= 16'sb000000_1010101011 && x < 16'sb000000_1101010101)  ? 16'sb000000_1001010000 : // m5 = 0.5782
                    (x >= 16'sb000000_1101010101 && x < 16'sb000001_0000000000)  ? 16'sb000000_1000010111 : // m6 = 0.5227
                    (x >= 16'sb000001_0000000000 && x < 16'sb000001_1110011010)       ? 16'sb000000_0110101110 : // m7 = 0.4204
                    (x >= 16'sb000001_1110011010 && x < 16'sb000010_110011001)    ? 16'sb000000_0101010000 : // m8 = 0.3277
                    (x >= 16'sb000010_110011001 && x < 16'sb000011_1011001101)    ? 16'sb000000_0100011101 : // m9 = 0.278
                    (x >= 16'sb000011_1011001101 && x <= 16'sb000100_1001100110)  ? 16'sb000000_0011111100 : // m10 =  0.2458
                    (x >= 16'sb000100_1001100110 && x < 16'sb000101_1000000000)  ? 16'sb000000_0011100100 : // m5 = 0.2227 
                    (x >= 16'sb000101_1000000000 && x < 16'sb000110_0110011010)  ? 16'sb000000_0011010010 : // m6 = 0.2051
                    (x >= 16'sb000110_0110011010 && x < 16'sb000111_0100110011)       ? 16'sb000000_0011000100 : // m7 = 0.1911
                    (x >= 16'sb000111_0100110011 && x < 16'sb001000_0011001101)    ? 16'sb000000_0010111000 : // m8 = 0.1796
                    (x >= 16'sb001000_0011001101 && x < 16'sb001001_0001100110)    ? 16'sb000000_0010101110 : // m9 = 0.17
                    (x >= 16'sb001001_0001100110 && x <= 16'sb001111_0000000000)  ? 16'sb000000_0010100110 : // m10 =  0.1618
                                                                                    16'd0 ;

    // Choose value of constant c based on input x value
    assign c16_w =  (x >= 16'sb000000_0000000000 && x < 16'sb000000_0010101011)  ? 16'sb000000_0000000000 : // c1 = 0
                    (x >= 16'sb000000_0010101011 && x < 16'sb000000_0101010101)  ? 16'sb000000_0011110101 : // c2 = 0.2391
                    (x >= 16'sb000000_0101010101 && x < 16'sb000000_1000000000)  ? 16'sb000000_0101000110 : // c3 = 0.3179
                    (x >= 16'sb000000_1000000000 && x <= 16'sb000000_1010101011) ? 16'sb000000_0110000100 : // c4 = 0.37895
                    (x >= 16'sb000000_1010101011 && x < 16'sb000000_1101010101)  ? 16'sb000000_0110111001 : // c5 = 0.431
                    (x >= 16'sb000000_1101010101 && x < 16'sb000001_0000000000)  ? 16'sb000000_0111101001 : // c6 = 0.4773
                    (x >= 16'sb000001_0000000000 && x < 16'sb000001_1110011010)       ? 16'sb000000_1001010010 : // c7 = 0.5796
                    (x >= 16'sb000001_1110011010 && x < 16'sb000010_110011001)    ? 16'sb000000_1100000110 : // c8 = 0.7558
                    (x >= 16'sb000010_110011001 && x < 16'sb000011_1011001101)    ? 16'sb000000_1110010100 : // m9 = 0.8949
                    (x >= 16'sb000011_1011001101 && x <= 16'sb000100_1001100110)  ? 16'sb000001_0000001110 : // c10 = 1.014
                    (x >= 16'sb000100_1001100110 && x < 16'sb000101_1000000000)  ? 16'sb000001_0001111011 : // c11 = 1.12 
                    (x >= 16'sb000101_1000000000 && x < 16'sb000110_0110011010)  ? 16'sb000001_0011011110 : // c12 = 1.2172
                    (x >= 16'sb000110_0110011010 && x < 16'sb000111_0100110011)       ? 16'sb000001_0100111010 : // c13 = 1.30676
                    (x >= 16'sb000111_0100110011 && x < 16'sb001000_0011001101)    ? 16'sb000001_0110010000 : // c14 = 1.391
                    (x >= 16'sb001000_0011001101 && x < 16'sb001001_0001100110)    ? 16'sb000001_0111100001 : // c15 = 1.4695
                    (x >= 16'sb001001_0001100110 && x <= 16'sb001111_0000000000)  ? 16'sb000001_1000101101 : // c16 = 1.5442
                                                                                    16'd0 ;
    
    // Assign value to wire
    assign y = y_reg ;
    assign mx32_w = mx32_reg ;
    assign mx16_w = mx16_reg ;
    
    // Counter for FSM
    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            cntr_sqrt <= 4'd0;  
        end else if (cntr_sqrt <= 4'd3 && sqrt_en) begin
            cntr_sqrt <= cntr_sqrt + 4'd1;
        end else begin
            cntr_sqrt <= 4'd0;      
        end
    end

    // calculate y = mx+c
    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            mx32_reg <= 32'sb0;  
        end else if (sqrt_en) begin
            if (cntr_sqrt == 0) begin
                m16_reg <= m16_w ;
                c16_reg <= c16_w ;
            end else if (cntr_sqrt == 1) begin
                mx32_reg <= m16_reg * x;   
            end else if (cntr_sqrt == 2) begin
                mx16_reg <= mx32_reg[25:10]; 
            end else if (cntr_sqrt == 3) begin
                y_reg <= mx16_reg + c16_reg;  
            end
        end else begin
            c16_reg <= c16_reg ;
            mx16_reg <= mx16_reg;
            y_reg <= y_reg ;    
        end
    end
    
endmodule

